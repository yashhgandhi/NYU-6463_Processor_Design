----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:10:46 11/27/2017 
-- Design Name: 
-- Module Name:    InstMem - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use work.RFPKG.all;
use work.DMEMPKG.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InstMem is
Port (  clr : in std_logic;
			addr : in  STD_LOGIC_VECTOR (31 downto 0);
         Instr : out  STD_LOGIC_VECTOR (31 downto 0));
end InstMem;

architecture Behavioral of InstMem is

type imem is array(0 to 516) of std_logic_vector(31 downto 0);
constant im: imem := imem'(
"00000000000000000000100000010000",
"00000000000000000001000000010000",
"00000100000011000000000000011001",
"00000100000011010000000000000000",
"00000100000011100000000000000011",
"00000100000011110000000000000000",
"00000100000100000000000001001101",
"00000100000100010000000000000000",
"00000100000010110000000000000000",
"00000100000010100000000000011100",
"00000100000111100000000000011100",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00011101011010010000000000000000",
"00000000001000100001100000010000",
"00000000011010010001100000010000",
"00110000000000000000000000110001",
"00000000000001000000100000010000",
"00100001011000010000000000000000",
"00000000001000100010100000010000",
"00011101010010000000000000000000",
"00000001000001010011000000010000",
"00001100101001010000000000011111",
"00000000000001101001000000010000",
"00000000000001011001100000010000",
"00110000000000000000000010011000",
"00000000000101010011100000010000",
"00000000000001110001000000010000",
"00100001010000100000000000000000",
"00101001100011010000000000001001",
"00000101101011010000000000000001",
"00000101011010110000000000000001",
"00101001110011110000000000001010",
"00000101111011110000000000000001",
"00000101010010100000000000000001",
"00101010001100000000000000010100",
"00000110001100010000000000000001",
"00110000000000000000000000001111",
"00000000000000000000000000000000",
"00000100000010110000000000000000",
"00000100000011010000000000000000",
"00110000000000000000000000100010",
"00000000000000000000000000000000",
"00000100000010100000000000011100",
"00000100000011110000000000000000",
"00110000000000000000000000100101",
"00000000000000000000000000000000",
"00000100000111011111111111111111",
"00010111101111010000000000011101",
"00000000011111011110100000010010",
"00011011101111010000000000011101",
"00010100011000110000000000000011",
"00000000011111010010000000010011",
"00110000000000000000000000010011",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000001110000000010000",
"00000100000011010000000000000000",
"00000100000011000000000000011001",
"00011100000000010000000000100001",
"00011100000000100000000000100010",
"00000100000010110000000000000000",
"00011101011010010000000000000000",
"00000000001010010000100000010000",
"00000101011010110000000000000001",
"00000101101011010000000000000001",
"00011101011010010000000000000000",
"00000000010010010001000000010000",
"00000000000000000000000000000000",
"00000100000111100000000001001111",
"00000000001000101101000000010011",
"00000000001000101101100000010010",
"00000011010110111011000000010001",
"00000000000101101001000000010000",
"00001100010111000000000000011111",
"00000000000111001001100000010000",
"00110000000000000000000010011000",
"00000000000101011011100000010000",
"00000101011010110000000000000001",
"00000101101011010000000000000001",
"00011101011010010000000000000000",
"00000010111010010000100000010000",
"00000000001000101101000000010011",
"00000000001000101101100000010010",
"00000011010110111100000000010001",
"00000000000110001001000000010000",
"00001100001111000000000000011111",
"00000000000111001001100000010000",
"00000100000111100000000001011100",
"00110000000000000000000010011000",
"00000000000101011100100000010000",
"00000101011010110000000000000001",
"00000101101011010000000000000001",
"00011101011010010000000000000000",
"00000011001010010001000000010000",
"00100000000000010000000000100100",
"00100000000000100000000000100101",
"00101001100011010000000000000011",
"00110000000000000000000001000111",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00011100000000010000000000100100",
"00011100000000100000000000100101",
"00000000000000001110000000010000",
"00000100000011000000000000000010",
"00000100000011010000000000011001",
"00000100000010110000000000011001",
"00000000000000000000000000000000",
"00011101011010010000000000000000",
"00000100000111100000000001110101",
"00000000010010010001000000010001",
"00000000000000101001000000010000",
"00001100001111000000000000011111",
"00000000000111001001100000010000",
"00110000000000000000000011011011",
"00000000000101011100100000010000",
"00000011001000011101000000010011",
"00000011001000011101100000010010",
"00000011010110111100000000010001",
"00000000000110000001000000010000",
"00001001101011010000000000000001",
"00001001011010110000000000000001",
"00011101011010010000000000000000",
"00000000001010010000100000010001",
"00000000000000011001000000010000",
"00001100010111000000000000011111",
"00000000000111001001100000010000",
"00000100000111100000000010000011",
"00110000000000000000000011011011",
"00000000000101011011100000010000",
"00000010111000101101000000010011",
"00000010111000101101100000010010",
"00000011010110111011000000010001",
"00000000000101100000100000010000",
"00101001100011010000000000000100",
"00001001101011010000000000000001",
"00001001011010110000000000000001",
"00110000000000000000000001101110",
"00000000000000000000000000000000",
"00001001011010110000000000000001",
"00011101011010010000000000000000",
"00000000010010010001000000010001",
"00001001011010110000000000000001",
"00011101011010010000000000000000",
"00000000001010010000100000010001",
"00100000000000010000000000100111",
"00100000000000100000000000101000",
"00110000000000000000001000000100",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000100000111011111111111111111",
"00000000000000001010000000010000",
"00101010100100110000000101011011",
"00000110100101000000000000000001",
"00101010100100110000000010000000",
"00000110100101000000000000000001",
"00101010100100110000000010000101",
"00000110100101000000000000000001",
"00101010100100110000000010001010",
"00000110100101000000000000000001",
"00101010100100110000000010001111",
"00000110100101000000000000000001",
"00101010100100110000000010010100",
"00000110100101000000000000000001",
"00101010100100110000000010011001",
"00000110100101000000000000000001",
"00101010100100110000000010011110",
"00000110100101000000000000000001",
"00101010100100110000000010100011",
"00000110100101000000000000000001",
"00101010100100110000000010101000",
"00000110100101000000000000000001",
"00101010100100110000000010101101",
"00000110100101000000000000000001",
"00101010100100110000000010110010",
"00000110100101000000000000000001",
"00101010100100110000000010110111",
"00000110100101000000000000000001",
"00101010100100110000000010111100",
"00000110100101000000000000000001",
"00101010100100110000000011000001",
"00000110100101000000000000000001",
"00101010100100110000000011000110",
"00000110100101000000000000000001",
"00101010100100110000000011001011",
"00000110100101000000000000000001",
"00101010100100110000000011010000",
"00000110100101000000000000000001",
"00101010100100110000000011010101",
"00000110100101000000000000000001",
"00101010100100110000000011011010",
"00000110100101000000000000000001",
"00101010100100110000000011011111",
"00000110100101000000000000000001",
"00101010100100110000000011100100",
"00000110100101000000000000000001",
"00101010100100110000000011101001",
"00000110100101000000000000000001",
"00101010100100110000000011101110",
"00000110100101000000000000000001",
"00101010100100110000000011110011",
"00000110100101000000000000000001",
"00101010100100110000000011111000",
"00000110100101000000000000000001",
"00101010100100110000000011111101",
"00000110100101000000000000000001",
"00101010100100110000000100000010",
"00000110100101000000000000000001",
"00101010100100110000000100000111",
"00000110100101000000000000000001",
"00101010100100110000000100001100",
"00000110100101000000000000000001",
"00101010100100110000000100010001",
"00000110100101000000000000000001",
"00101010100100110000000100010110",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000100000111011111111111111111",
"00000000000000001010000000010000",
"00101010100100110000000100011000",
"00000110100101000000000000000001",
"00101010100100110000000100001111",
"00000110100101000000000000000001",
"00101010100100110000000100000110",
"00000110100101000000000000000001",
"00101010100100110000000011111101",
"00000110100101000000000000000001",
"00101010100100110000000011110100",
"00000110100101000000000000000001",
"00101010100100110000000011101011",
"00000110100101000000000000000001",
"00101010100100110000000011100010",
"00000110100101000000000000000001",
"00101010100100110000000011011001",
"00000110100101000000000000000001",
"00101010100100110000000011010000",
"00000110100101000000000000000001",
"00101010100100110000000011000111",
"00000110100101000000000000000001",
"00101010100100110000000010111110",
"00000110100101000000000000000001",
"00101010100100110000000010110101",
"00000110100101000000000000000001",
"00101010100100110000000010101100",
"00000110100101000000000000000001",
"00101010100100110000000010100011",
"00000110100101000000000000000001",
"00101010100100110000000010011010",
"00000110100101000000000000000001",
"00101010100100110000000010010001",
"00000110100101000000000000000001",
"00101010100100110000000010001000",
"00000110100101000000000000000001",
"00101010100100110000000001111111",
"00000110100101000000000000000001",
"00101010100100110000000001110110",
"00000110100101000000000000000001",
"00101010100100110000000001101101",
"00000110100101000000000000000001",
"00101010100100110000000001100100",
"00000110100101000000000000000001",
"00101010100100110000000001011011",
"00000110100101000000000000000001",
"00101010100100110000000001010010",
"00000110100101000000000000000001",
"00101010100100110000000001001001",
"00000110100101000000000000000001",
"00101010100100110000000001000000",
"00000110100101000000000000000001",
"00101010100100110000000000110111",
"00000110100101000000000000000001",
"00101010100100110000000000101110",
"00000110100101000000000000000001",
"00101010100100110000000000100101",
"00000110100101000000000000000001",
"00101010100100110000000000011100",
"00000110100101000000000000000001",
"00101010100100110000000000010011",
"00000110100101000000000000000001",
"00101010100100110000000000001010",
"00000110100101000000000000000001",
"00101010100100110000000000000001",
"00000000000000000000000000000000",
"00010111101111010000000000011111",
"00000010010111011110100000010010",
"00011011101111010000000000011111",
"00010110010100100000000000000001",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000011110",
"00000010010111011110100000010010",
"00011011101111010000000000011110",
"00010110010100100000000000000010",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000011101",
"00000010010111011110100000010010",
"00011011101111010000000000011101",
"00010110010100100000000000000011",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000011100",
"00000010010111011110100000010010",
"00011011101111010000000000011100",
"00010110010100100000000000000100",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000011011",
"00000010010111011110100000010010",
"00011011101111010000000000011011",
"00010110010100100000000000000101",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000011010",
"00000010010111011110100000010010",
"00011011101111010000000000011010",
"00010110010100100000000000000110",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000011001",
"00000010010111011110100000010010",
"00011011101111010000000000011001",
"00010110010100100000000000000111",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000011000",
"00000010010111011110100000010010",
"00011011101111010000000000011000",
"00010110010100100000000000001000",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000010111",
"00000010010111011110100000010010",
"00011011101111010000000000010111",
"00010110010100100000000000001001",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000010110",
"00000010010111011110100000010010",
"00011011101111010000000000010110",
"00010110010100100000000000001010",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000010101",
"00000010010111011110100000010010",
"00011011101111010000000000010101",
"00010110010100100000000000001011",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000010100",
"00000010010111011110100000010010",
"00011011101111010000000000010100",
"00010110010100100000000000001100",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000010011",
"00000010010111011110100000010010",
"00011011101111010000000000010011",
"00010110010100100000000000001101",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000010010",
"00000010010111011110100000010010",
"00011011101111010000000000010010",
"00010110010100100000000000001110",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000010001",
"00000010010111011110100000010010",
"00011011101111010000000000010001",
"00010110010100100000000000001111",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000010000",
"00000010010111011110100000010010",
"00011011101111010000000000010000",
"00010110010100100000000000010000",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000001111",
"00000010010111011110100000010010",
"00011011101111010000000000001111",
"00010110010100100000000000010001",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000001110",
"00000010010111011110100000010010",
"00011011101111010000000000001110",
"00010110010100100000000000010010",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000001101",
"00000010010111011110100000010010",
"00011011101111010000000000001101",
"00010110010100100000000000010011",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000001100",
"00000010010111011110100000010010",
"00011011101111010000000000001100",
"00010110010100100000000000010100",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000001011",
"00000010010111011110100000010010",
"00011011101111010000000000001011",
"00010110010100100000000000010101",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000001010",
"00000010010111011110100000010010",
"00011011101111010000000000001010",
"00010110010100100000000000010110",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000001001",
"00000010010111011110100000010010",
"00011011101111010000000000001001",
"00010110010100100000000000010111",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000001000",
"00000010010111011110100000010010",
"00011011101111010000000000001000",
"00010110010100100000000000011000",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000000111",
"00000010010111011110100000010010",
"00011011101111010000000000000111",
"00010110010100100000000000011001",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000000110",
"00000010010111011110100000010010",
"00011011101111010000000000000110",
"00010110010100100000000000011010",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000000101",
"00000010010111011110100000010010",
"00011011101111010000000000000101",
"00010110010100100000000000011011",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000000100",
"00000010010111011110100000010010",
"00011011101111010000000000000100",
"00010110010100100000000000011100",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000000011",
"00000010010111011110100000010010",
"00011011101111010000000000000011",
"00010110010100100000000000011101",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000000010",
"00000010010111011110100000010010",
"00011011101111010000000000000010",
"00010110010100100000000000011110",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00010111101111010000000000000001",
"00000010010111011110100000010010",
"00011011101111010000000000000001",
"00010110010100100000000000011111",
"00000010010111011010100000010011",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00000000000100101010100000010000",
"00110000000000000000000111111001",
"00000000000000000000000000000000",
"00000100000111110000000000011100",
"00101011110111111111111000100001",
"00000100000111110000000001001111",
"00101011110111111111111001010010",
"00000100000111110000000001011100",
"00101011110111111111111001011101",
"00000100000111110000000001110101",
"00101011110111111111111001110100",
"00000100000111110000000010000011",
"00101011110111111111111010000000",
"00000000000000000000000000000000",
"11111100000000000000000000000000");
								 
begin

process(clr,addr)
begin
if(clr='1')then
	instr <= im(0);
else
	 instr <= im(conv_integer(addr));
end if;

end process;


end Behavioral;

