----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:32:21 11/27/2017 
-- Design Name: 
-- Module Name:    DataMem - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use work.RFPKG.all;
use work.DMEMPKG.all;
--use ieee.numeric_STD.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DataMem is
Port (clk : in  STD_LOGIC;
		clr : in  STD_LOGIC;
		addr : in  STD_LOGIC_VECTOR (31 downto 0);		-- This is the ALUResult
		DMIn : in  STD_LOGIC_VECTOR (31 downto 0);		-- This is rt_data from Register File
		DMOut : out  STD_LOGIC_VECTOR (31 downto 0);
		sel_wr : in  STD_LOGIC;		
		sel_rd : in  STD_LOGIC;
		l_arr : in STD_LOGIC_VECTOR (127 downto 0);
		din : in STD_LOGIC_VECTOR (63 downto 0);
		data_mem: out DMEM
		);
end DataMem;

architecture Behavioral of DataMem is
--TYPE ram IS ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
--signal mem : ram := ram'(x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000",
--								x"00000000", x"00000000",x"00000000",x"00000000", x"00000000", x"00000000", x"00000000", x"00000000");

signal mem : DMEM := DMEM'(
"10110111111000010101000101100011",
"01010110000110001100101100011100",
"11110100010100000100010011010101",
"10010010100001111011111010001110",
"00110000101111110011100001000111",
"11001110111101101011001000000000",
"01101101001011100010101110111001",
"00001011011001011010010101110010",
"10101001100111010001111100101011",
"01000111110101001001100011100100",
"11100110000011000001001010011101",
"10000100010000111000110001010110",
"00100010011110110000011000001111",
"11000000101100100111111111001000",
"01011110111010011111100110000001",
"11111101001000010111001100111010",
"10011011010110001110110011110011",
"00111001100100000110011010101100",
"11010111110001111110000001100101",
"01110101111111110101101000011110",
"00010100001101101101001111010111",
"10110010011011100100110110010000",
"01010000101001011100011101001001",
"11101110110111010100000100000010",
"10001101000101001011101010111011",
"00101011010011000011010001110100",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",--
"00000000000000000000000000000000",--
"00000000000000000000000000000000",--
"00000000000000000000000000000000",--
"00000000000000000000000000000000",
"00000000000000000000000000000000",--
"00000000000000000000000000000000",--
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000");

								
--signal memaddr : std_logic_vector(31 downto 0);

begin

--Store 
process(clk, clr, sel_wr, addr, DMIn)
begin
if(clk'event and clk = '0') then
	if(clr = '1') then
		mem(40) <= l_arr(127 downto 96);
		mem(41) <= l_arr(95 downto 64);
		mem(42) <= l_arr(63 downto 32);
		mem(43) <= l_arr(31 downto 0);
		mem(50) <= din(63 downto 32);
		mem(51) <= din(31 downto 0);
	end if;
		if(sel_wr = '1') then
			mem(conv_integer(addr)) <= DMIn;
		end if;	
end if;
end process;

--Load
process(clk, clr, sel_rd, addr, mem)
begin
--if(clk'event and clk = '0') then
if (clr = '1') then
	DMOut <= x"00000000";
else
	if (sel_rd = '1') then
		--memaddr <=(to_unsigned(addr));
		DMOut <= mem(conv_integer(unsigned(addr(6 downto 0))));		--DMOut <= x"00000010";
	end if;
--end if;
end if;
data_mem <= mem;
end process;

end Behavioral;

